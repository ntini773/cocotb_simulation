module simple_dut(
    input clk,rst,
    output op
    );
endmodule:simple_dut